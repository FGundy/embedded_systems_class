----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/10/2025 04:12:38 PM
-- Design Name: 
-- Module Name: hw2_question3_selectedsignal - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity hw2_question3_selectedsignal is
--  Port ( );
end hw2_question3_selectedsignal;

architecture Behavioral of hw2_question3_selectedsignal is

begin


end Behavioral;
